../sw/rom.vh